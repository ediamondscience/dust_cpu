library ieee;

package ram_loader is
    impure function ram_load_from_file(
        load_file : in 
    )
end package ram_loader;
